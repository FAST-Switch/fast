��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��� o�tL��nàZ�mv6�9��g�q���V��wy�Vi�f��:l*�K��ņ2'x��BG���da�l�A��{2�������Fa��P�(V�qF� �:\%u�f�WCy��VQ$-;t�EA�A�K����M�#�b�<��$hW}�_v�G�1��1�"����K�1�A}#|CU�Vl��gm6ڜr�C7��L�n�;��$yB��)׬j�9H�7w�����,��%���\D�@��d�BY�������LZ%w���%kG�t��j�;<W��������Y�g�����Ɨ<%N��'$e�h��h��8�qoQ�4]�A/Jz�!a;,�%��$b ��?��!������/3� �4�y�z�u.���#��ʭ�+��u� ���Z�T���84Z�	���8���sA���v�Sߨ�#t�y�[�p�ˢM^��r������EV��N�̼81��$,k��vu^T��[��|9ܷk��3���қH�H�����ɷ���R�r +�����ʮ���� <�j�$� �%�[�f?��t���N��Y�tʈ-�@��tk���j�9�m�8�u���ٺ./�W�ҒՈ�[ur���i{<���艚��D�����W�s��|�Yz�a<<u啥|�+�'�a�q����|�x[���iߌ�����q�H��S�# ��QK�\�:2���x1>8c(C$ܪ��Rɽo�$�Qo��=[�O5���?���RMj���f>�Ǆ��pd�C�8,0~H��b H���1Z�Ϗ�R.�2���d��ۊ\�����>јA�r?�y̴�,�\o�:4	��M��C�ڰ5\P�y^��d�F/� �_�]z��=6Lw ��)��U�8>���<m�`ϔ��|WvXr1qG��q��Q�])�@��a�����	a[9�	��E�|��}4��Ŵ��~��.������~��ڊP��:6�n]���~9��؁I:�{�h���I�a�7�5ЅJ[1�M�L�.(���&��(��U1� "j� ��o��g��r��?����=X�Rm�Uk����B����B�L��U�0r�����t�=���%���SoHehBL�kv7S����£��A�+i�u���]F����
k��<A~�C���������*�xq�.�8�N"h�}�����p*p�c�XQ�_B�'ɓ�<���o9�s�TiI�IP7t�9�/�f�f�&i@���&�r�v���V�b�rS�X�\�5�&�^��j����zH��)�i��}nfv5�A�n"u���Zh�e�R����Ԅz{h��~�\l��|�P��(D�I~�A��n��}V�|��7�I�hl�Q�q&5S���k�!ִyN:|�{���Q�� �1�d@�$l����s����M
K�<�>�$�Ȫ ���6�q��F�353A�b�[�"Q�uC�s��8`�vY�$G�L��Ul�`B�4�I��Y���(p�v�c���D�N�޵��x�I�;"�b��m���=��1�qa* ��dy�6��x;V�m`zh�e�>�j�+!0)몴��tӻ�{�U�`ʱb�k��#� ޷͟9w=�vX'�Cı�"2L�`��&|�8B<Z���U�#M���*���zX;�s���{���*c���{?��)�;X�* �|�Y]G��)
��Yڬ�����	Ws�:�&��@J3���p����S��t���HzI	����	�<�{]��t��7}�lm=��Q�Ƨ>�r���[,^��y?��F�ش����.�는K_X3Vb��ҤH���d����@�%�2�Q!����l�d(�p�XФ��d� �K0�*�G�2aK���Dl���G��7AA^#W�`��Q��r=&�pI/�|J ��;*7\w�lxi���e�S�FO�f��E��C�ܐC���#�dK��)�]b'AT&�nV��ZV�������A�!nt�Ja(eQ��)��(�AQ��ߋX����>��rQ���N��\�ь�1�������C���^��� ��J�ƹ��g�T-Ġ�f���Zº'w�;*��"U��75��@4@u����A���it�lM�0d����b�G=�C���ە�'�l?���&� ����7�&l(�ಙ����_5�\�|{�:��3\b��s���L ���5q�v�0�Nh��N�A�w'��Åymr� �8�� ��<������5-�m�?t�^�HMX#����a�����TlӤ� |��;�iM}Q)VH1}��O
6į��X��HTO�Α��%c� #��7����5��,!6ͧ���|��]P�����!�e�n�M�@;-&�Y{m.��͜&�듖�g��z3j���p=})N�z	R��T���:����m��#s>�^����(s��}�pUu�3�٥K���� ش�u�$oa_�E��q��/4�����W�W����4	���4��ch�[Y!� °�#���1�9'xҞ3�-�!Ru*�M�SC��3�+(����鵸��1r����?ymP�΅���ljm��
c3��x���Y9��Å?�3�i���E���A����ֺE����tF��J�?nJ�zY����I��>���8ė�(�����s�si��
 J�w��2�����XK���}EFaJ�5���"���Re9S��ʤue�Z֭x�-�n�pyC����G�u�Ι�G�P�d��s�� ��3QW�X���6bT��"�� Uu���kT����m������C/���Hh�|]�K���Ly�wSs�|��Ƞ}J*��Z}P��&��D�)F���I�^��2�싙�v��?�l�DV���9�?ő�����a;��K7��ꢯ������-=Ng��A��\�)���-�XB��l5	�T�t<�q����^��Q�}�s2sF_Mo��ŗ�Y�Lo����_��+0���ӯ�ә\�;d��tR���t�J+i��t�?0>�x.V���!".�N��z��st��Q�H���d��~A8hQx���"�z�Z<�m�Ha�ۜ(J�vEsy�Nbɘ�`q�l��څ�O#X��/��y}P	 ���Q�ZE�.x�b��g��5�[�U�b���e��3}cM}6���O�6�9�1 �&�.x�!�y��AU����������Ի�ſ�l[���":��,�v���`�ì��@|~����3#����`5��Rj��'���hu[u�_�J�'�r����L��ϷvA�ܘ721���Ӂ���Z� �+ݱZk3]��SϚ�o�n�nG�ّ�zc*BŪ/Lh���&��!u�]n�~ o�6	q4as}��
�9޾�p\4OSc�U5�4��&j�&�g(׊(ƧPQ^��YhlCUI�s�����!��ȇ;�P٣7��E�����nkKѸ-�O��Fr/�k���H� �����QACv���/����QY�3�N�#@�b*Κ|���r�P�:��G~��P�j���5=f��8ƕ�^�Ų}�Hlðǃ���  L���Ώ~�0���������@���H]�}���k+�}�~����ue���^Jlh{h&p�>�,�7rN��&�=n�N�D�L�(�Co�sN�/�����q���i�����E�h�+�B����$ѱ�����Q���x�-�+��	�Sgx�=P!*�됀��ܜMcrs�W���fS2ā�9�?A�U|�d,R�����Fs;��^ї4��O�gc�j{>�Ɠ���ʅX0����SU/z����j�K��	�ȩ��K�Fbdj.��Gl��)R��;M�r�YK.��$%�΁j�JP��8W�I�{�@��>m����6ج[��������'V��h2��&��G�����?��(�����
g�=2L�i�f��ٮࣶ�a6uYn/~����0j��A�ZC>��z�eW�T\�@~�al5Ô|'\ޒ`+d���}؃���Е&)�J ��ņ�Hȇ^BF|
-r弶��u�M���/,���o��6u�w������2�%�C��i����X���A���:0�(9�]��j��c���l{3 &/hV�x��S�B2�y��+������������1�D#ͮ�,� ��/Q7�@��'�ݽ�wZ�ޕۼ����c]4u���|�x��O���fO⽯��