��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?�T�RH��'3�g��	o���:$$LEχ�K���6k����8��>����Vlˡ���s��Uޯ��	c���D�?)��#�@W�{; ���͐/���O)C}�C�>�؁eΕ�Y�8�ﳻ��/N��;�Kw�O�h���+�5uO c�7w�X�8�VĪ6����;�!jA:I��{�dD��Z�T%��"*�!gǽ��阬�ϋgԁ�zp���"�2O�w��qݣr}��݄�x����e�RʿH=҂
����?	(I��7D��a������o��M��룍L�ةx,�������4��_�h���wa�������"\�9E�P=�����'a�ZѠ�ٞ���!�V�)L�AΛ�׊n�jRR�(��:��@�ny̰T8A��L=�OD���yE���澒�7�lR��R�
�6Hb��������9'Gu�=�����D?|�v�#%�n�C���5�����6rk�	�Vc�kC,�"�8a�Y�R�y�@B|�N�ʛ`�XL<���r��He�����±�+	���'�[q�������nȝ�TU_�����b��ڐ��|��KT2��K�uߵ���ۙ�墍�T�����p6Ҹ̹���i�dҜC�cE�2n�]t�YJ�e���+��ddO�t���`QI�8�$D�t�=�܎*Ï����[�H1'5�o:����x�<�d���Ms�v�3��5P��[M�ҏ��3�yc98�������giT~�gBN^�+@�������f��R�@�1�1��r�p��G��1�~d�#��վ�m���YSʫ-���䱂���RA{L?̆�UR�����!6B�ѯ�w$����v�����D�!K�1��q��~��ǆ��O]��ɏ$i�[��w��$C۳��y���]� ��c�v�r��5�|�jY�(]�3�ՙ9�Q�5���1��6t�����m���^ň���iTh���7�+� �V���^���]y7�֯���Y���]���"UVd�5]�l����6��R�J[,���ɺ|c�C��Ñ��wc�����J+/���q�Gd�����.�OW��
)?�Ո��(}V�)���ʠ�M��f�<x�Q�T��i	�}��X���c:��R��$��&5�5sW3"����o�_JM �[�ւ��qx|�=x�4�O�z��4?zd��;�g]�?q�]i�#�H��B�/��!�J�G�rk���RM�Tn����<�k�b{n7³�nm~��v�L��{���F�����AE����sLԑz��̓A�X D��������^�q�����Z����knP$�j���Z��ni������q�*9|}2�猁�~@�Ou�#J�5=��:+�s\+"�펂�'�����rϦ�&\���\�.�|�`�I&Púz��9���O��׻��%ś��� H��,ƾL�<"�.+*��X%�/L�\鱰��	%:}E��^3uSeW{���m�7��'���q�?Z�Hk��Ñ�$��~�EQ�����./ԓ�Qg�A�(���#�������J�Ǌ�ؤ���Y�N�oNν��!i !LU� h&�	J����pS/t����iϔ�\y۽z��.��ߏ�#C�����7V3��1�d����� �юr�/:��m���T�0%�i��oQ=�27ՌL�T;��yc�p��{��9���8W���Y��~�6��+T�m:DD�����<���OV3��*��D��6c�uЍj<J��AM �7R.�$/�k^8)�_&(�� ����u�aM�X�<%z����Iܷ%�pn��"��+X�ZF�ň�UN�&I��Gmp^ؒy��^�U�o���hK�m�A+	j��7=��t�v�S�H����G�%r� �3���b�����aͤ]��V�EYX�$���������({tY�l�DƳ┺�60��+Q�t�5^򻌨K�9'
 $��*2��i"֗Z��lɖ�2M}�)��59�)�6�� e��( h�i.�f�ɒ�L�״Gte��"�qV����(��a3�p ���2I�é���d��՚�V�^��ߦ�?)tЪ!�B��R{�1��@vk˯�Ut���M�8�j�*�[�Z���b���ꪺ�+�"d���X�c
�]��ġ�ͯ�= s�:����I����Cw��ð��K��cd��g�Vn�:�&pH�?\��Cc��~@1YC�D�Y� s��9��&2��ߜ�t����N}5�C�Hu��l�ư�J�]e�՗{9���uҘ-.a����-�(C��X��C����8�u?�h��t��oK�:W�"��{�W�m�=m���v��Xv��.�­��*L���^c
�*���Y���8�JC�`�A;�Æ��欶O�kn�YO��
���U�=j�uf�Ҋ��f�6b�q�w����k��!Ş���w2��W9+˝Ш0Y%��|�h�l
�.P�����-����UD������<0�h :,���M�b*�mwZ��xrZ�q1����e�\����-�
�5�:�@�U`w�;!��2�L�wt7��6<<�CžS��똩��]&�T������!J��ARL𩂞M�������/���k��WӘS��4�6q
"Eb�� �X@9�o�f!!��YN��E.E�J�e�	�?*{H9WŰ�Q���QL|}~́	"��'�*�0Z��!�P(w�[�����;��tUfK�.�}���"�W�=?�"�����s���d�P��ʂ���K��6�[� ��>����}|��~�N���=׏5����xD��tJ����,ꍗY����a�˾YG��K�� i!Q �G�я�*8j��!o[��a�������|&mr�J�Y�-�z�~�xaT��s��]4 �G�9�*�`��z�˜N޺� {�MJ'���R��#Y�@�b�4�FZ��J�~K��6-0oS�du���Oκ��h����U�sޛA��9�K	+���	�w��Q ���X��h-RiL8:�{�[�^'�w�c�K�'f��4��i�N�v��#N�a8 �q~\��O悮/��.S*$l�[��S*1��M9Ir��NQv:� �h^
�	��఼��/��ՠ	�����;$���]�I<��n��}���Kc~@���E���N�T��a�󢐒���3�}\��tr����V��aO	s��n��V��&��w
&�<k�OD������E��S確�1�1�έT�v�7�P! ��n���D���}�����zIN�ߖ@�K��R�q,���L���K�!5q�:M�.q��ޠƪ���p!G��ݏ�/h�ye#�&�LeЦE$��A��DS�6d�ӝ2Y�l�o��'y(A�<�$��f%�b�>Z�}��w���QԸ�A��Ɏ�h���<t�d�MH��}�:a� XZ�>͹]})�UtJƵ\���S��&�ЩW"���A]�������ih1���4�iᖟ{��y�������
����Z�k��xG�5	[1z	�uD��i�o��D>�D'8e@�7]��q/��%�y�b���ؐ��J������@��d�����ư�b���{�r-��4�5�w4F��2��@��ԝ.���>ƨ7�(�b�mVΕXy�vOo>�Wە��{�MKf@|�Oq4�Y�g���H��}��z��P\颍"����/ ��k(yRLU�� h�x� p��J:�����.=�9���f�#ӕ�邗J�+�����޽��6�����<�ݹw����|@蝺 9邅�we����s��N<d��x�v^
�DП�r%� -�0�_��fU�_���{��<����)�Dm3A̺���9Ƨwۥ�'
��,�����.@�f�|J�w�%��k��}�O*u��(f�/�@Nۂj�(��23�^P�v�Ή�9iӎ̃��$��yu��ۋ���M$6����~)��ϟ^V�;l��s��,ܴ�ǘ�,��i�?����ҁ���3H	!��V���	q�vp��)�6����EDZ.��;�Nn����`�ی���S�v(F����aӦv<�7�cETqp���	���D����ٙ�_8N�o)γQ�MC[�/]��~$:f#tD�1@����'x�>8X����v���,�'��vc���-��:���UWDy��I�Ū����/-p��q���I[)_����=��+��+`
Ьv,�;��_�F�ӈ�����7ɰ
eܱ�e{��5���