��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D���3�'��aE��
�<P���ӹ�`^�dfFVN��l�Z�	��Xkɑ<�|���X@�=A��4�w��a���F�B��^E%?��}����(�d�8�z�-(��Q� ���Ps�Y�Xg:�y��7h�!Ϯ�����F��5c��J��q.�Gba��8W	)
��l@zB�P��L�E3f��4�5ޟ�jS��{_�e��ќF���#m`���WTÿ��x��3H�ovd&Ź`M�"���<�U#�� ���[��z%d�}��x(�<��Z�����F_�V���k3�2�����J,Z�Dj��A�#�6z2�����l��}��8S�<N�į�����_(�?^�q��7R�r~
4��ee��u=��J�gbA�%4F�>6��5֠T��٥��	�8����>�4n�|c�C�W���0r1�O29ظ�Mwtv�`�N~ �_�Xr�,�yX�U�R��\���}yg��P�l4�~ߙ���K̅�?p�p)�`t�:�'Ȓ�
�:&�u�K����ʥ���=�����ણO�~#r�<�{lAP��2UM~G��f�,�k�#Q�;���Lm��gt���څs^C�L`�p��g)�÷�&-�K␕c�?d
-K9���Z�܁a�y�p�4�Em�ǘ���� � cb��b˹>c����������&L��UE��)΅V!!�� b�{�����J:-�����!��ei�.�	��!lCq��w�k7q}���:�.�i�_�}P~)$�G��_1L ��ۆOOS�3��ӗ���?�T�RH��'3�g��	�	��U��b$�n�JT�3 X���w�ܶ�42A#0�Y	K<�+0� K-g�����घ��A�d�N�oj6�H����:�qc4���u[�-���Ht�qC�m�]x�l�{��� �@�0e�[��������wG�Fď���X��fT���MW��I]Bo��a��R3�z>8$V#�|<KQo�FM��_V#�nƤfTL1p.��7/-�/���+���Q �Q�G�=�I�p�T��}2E�'ff��@x�r��ޱ[6^�\\ %�i��u��Y!�����*�p�������s�g�m�d�Xs�p(�]+�8;swvx˻-�⧃|��5t�D�L~�~�5�5�W��![y�:	r�[I���_��Pq� �G-r{�{\�x��&f���f�a<�-���Y����Q'��t�A�:W�R1y�j��Jr��
�vE1{��o��ŧ�|� ��Z7���~21�ȫa��.��c[��f�# uQ������)y�����æ���F�����UhOS�33�-����UP^xY��hB����g���p��H`�"�Q;�cι6��׋X]�kh�^�;2E��_SP���߇������=�B�jf%:�Ӡ�0I�6��˸U��Ơh��7& خ��3���\�&t4��4~@����[�4�{B��^])�&�f\Ԥ� �� $F���@����.�	���f���@�5�.$7���%���g��mk/"���5�{�9b'���.����������cH��B�*6��Ds�}����9���Wfz�����öh�d��_2Ql��<eZx����Zʲ�(��q��dú�����c=�E@
��BG�͜�u�v��I(@���t��=���]�U-�~�BA����O9b� ���eϳٟv)XӶc�ҘQ�xC���G��-$�ẜ�>�.�;`9����r�5�)���E�������_��
��x[b�
˫n7m��<>�a�kp�7��.�WIX!MK���@�5`�h��-zG��{��Ӽ�� �9���������-��U ҋ��La��6}uAW?I�xL�/����Gi�u1Ou����ې:uV���c1���m\�ppb.�B�����nP&Dh0{��dfz�nۧ���r�V�����;��\��[�3��)Df%�V#]?�������a Vjx�~��c�1�/�֥|mŋ։Z��my��ꩺy}v�/%�O,m<Bc������L��90���9�3�<n�@q�n6c�qTc�Lk��)i����Z�*�t��[h1>8�6��h���g�e��@,פ����O���*�$�B�@�DJ�_E��K^�g���9�8-�R�d���Ⅲ��+Ֆ��r����l�o��V������i��н�/���lׄ�و��4���?��d֑��Wy��7�s�rP�`_gh���z����xUJgP���b���Z J7%��2K��$�~�G�V��*@B[���J�������3�R��%~����ol���d�=�$DB��B����BbP>�C�l��F]EK�^�x��10��RY��N��,3E2�DB�Ti,۟���OL�^Ejz�
�yn=umLY� e"��S����6�x���|�v���+���ʢ`�5M)֩L�S:"���Ϫ͍��=�Lڷ����t(���|#�-G�
�����A���,�̋��-b���2��9>�]�F���7�W�cIƧ�_�3�ͪ�[={pt7b�NPn��Y�g��Z@�_ɋ�r�}r0Χ�xn��^�g$ƻn��������w߽R��\�oe�aw�w�dr�	%�#�Q�4�����O�8J(5Դ��"�m�VƦ_��ˠ<Y`cvӥ�С�~Ļ|!�7?�"_�m��C��m��.Sp�[�^���1�s���W���P� /	�V���J��$zE�l���)g ��l��q��@o�$kjȳy�� �%�[��@�w�6�Q�/�9,�OBmR�EV���P�M���c73�wI�'��D�nU�<�"�����s6h��A�ԽBogi��k���9�Gn�+ǫ���/�U�x��
g'Vtu³���~r����d�E;�5ۍ���N�?]pOKVE=������t�����=�T���o�4��O�nk�0r&}2(�Xn]3`Aف[= ����D�� l��E0����ޭ�d��b���A��a��oP��G�"�0m2��7���O��_�$1�������wӊ�]M�p2�9\��IO!��V54������.�)'�<�N�鹗̬חy
#v���ttT<��7��c�8���+�\�a�b]r��]�0��	T9����+��椱*i�mo�h�.��@\�9�C���P`@��I�"-?��|(�k�u����)׏����_ݸˢO��N����	�ٌ�\�>�<��	/N�GhJ�hװ��CA�`��Z�
��(n��àe�ţ�r�m��@(z�-�z+�����3#�u/��VŪ�ؓ��[����=��r2��P�ը�23��`��������������Y���yД��-P���։���Zj�bZ����6�3K��l��=�:hD\#v!��/��~��B И���J:M��f���~s��>�n.m�$H����O� #�J�GO:9�Q�^X}'a"f��2}N��R����#��Ş]��/��_E��N� ���-@3�J9p9�	o��
�".�C���b{�ԝ,2&��4����b���΀	N�	Z�$d�>���6Kk/��M��OX�n?�3���|���NҜ� ��P�%�s��˳=,�o��_��߭�.$P�m�C@�|�t�5^�����`V�p�ǵ/bI���koZ�B���q�4V���ǻ����ԗ�D\�A�{V��䩍n�=ܨ���,��%������]�.G�T���7�b�����>^̑� ��1���	#۽�b�`1���Z�igߡ��gr��9b�a.C�/����i�'���?R�P��:>p�6,<�w��������<�����h�gᶠ�JE=e�:�a�%��d��Ք�\Lrn--B�{�4��l}H�����M�|݇]�j���^��1Yf��*9���uJ�m�2�5�W7<7�9�3I���Q�j�Q��'c���R��M�V����Fr�s-�v��2�'\ho�J���u{�:W�=�s��W�њ��W���0cxޛZ�/6�����_�%�A�aӓ�2/�dн����o~�u��������Յ��P�ʄu�z2��*7S�������� 'k@Άh��a��%u)���Xi9ĺƭ}V��5ؔl[���~��?B������A�n'�ؒz�_NL�S�{O��=�˶e��G�ܻ�2�T�ā$��J-��+��Ap.�r���T8����up2-q�&B�U|�O����I���-�bK�d���jޙ�2n����1b-Ah�C�z_�  �{M��\<�����:�hy����P�T[��(Q�����s�ᗐ�B1]�]G�6eH�:� 0�S��pOI ;
��!�O<^���2������`�	�`�Y�q�"��rjd��i��0ջ�❐�} �Q3��ռem;�� ۻ�E6{�}�I�Y��.��G+J��0��U��#Pr��V��+�"
�1�w1����.
�ҭt1<���=�;��j��9+e����$�*`!<�5�Q<�ٗu��z�����.μBa�)ʼs�>ӵ^�Ӟ\�3���&duE77�W��3]�ԣZF�}%̪>!p�v�,���ū��F��N�O��"2vj�d��-�ۊȭ dR�+K$��C�/C� $����
�tcT�v,���j��Ty�q `NH<��M�D󥶺;��/J��I#�5�m�-��k1P9���}j�2���B)���TBvQ`�.	��������f��)�$I˟3��%��v�#�lW���=�{��0���L|���Zj^�MEc�|�\�J��E��U8%��u7�>���)�^YY+ fވG��i��b2��c���ோ��v�Q]��VT���]��hsJ��)������n�	���q>B)9��"͔� ���[��v.�/�!�:CV	�^�G#��B���J=Y]��Gm/'���Nx������9��E%�̨G(��D�71n$�1�s��Z�*��f��N�P��hCF�}N�\��^y��+%o��t��üYx�w�CJ�L�!!�GȌ���Ӥ�h8��G��-��f��G�)�F��~���
��OA ��q|@\�ʄ8jJT|����im$܊Aæ�X<�o�1�Ơ��Z����DKڈ��_�}4d��\#F�4���mez	N��Ua7�
s ��x�����U�vS��Pܫ�Y�6# �ل�e�_{�d�J��r4"�E��-Ax��L΢�$�J�b#4e�T:��T�����)�� �<�����cwf��6��*ͱz�E��ȯn����d�A���LBJ*A�ͽH��yvFs���L��@%�QIK:Q0,r�����g6���ߔ��Z�C��.|HU`FZ�������\nMqO�scP��,�	Ҭ����y�w��I�?��G����F�Fp�\�z�ԿW�$)*�0����~E�|�l��� 9V�@%/���U:�L���+%���}�;:B%�g}rc��r���Ȼ[?ٖ�/L�:tC.|z�S�!��ouZ�gc�š13���r�8惷LlZj�o��0�lb29��ǎ�h����,U�^�2���sucx�}noc
`0E��Ѫ4��p���N*ߍ��\�ش5���,�Ht��O,���Y#�Y�\� 3�
u��o�	J�	8��@Y`���q�lq{�G'z���X���KH��$�O<���Uˈ@&���G��<��f4d��!\c�� (`�����Ӻ�~�lYk��uT���5��σ�$D���;�{�z����n	�Y��3_I�y9%�[c�&�q������u5�bI�V��4P����q���(!s���1��MJXN激]ہ+-�ᬫ����>:�� u�*�x����m�Gv����U��}v��G|���Cnz�4k��w��/H����2��۾*�j�%���]�7 �oS� GD��ڃ���2�qS�q�c���%�_pL�`���Ni�c�G���t3V?ߩ_(�3��L]�O{�m�暯�~��㒑�I
qO�m�ڋ���{���B�1���v�+6��z��4���E�m�R��v��<�M��-�:�w�#�*k� -�2��Hǁ1����.�G�chh¦B�OQr�������=B�O�a����=y��=Ǌt�.z���Ŵ*�N�s��� f�V����Oc�M�V����S_��g��7�s"�3�����������M[>�~>="�����K;s�6Χ�I�"t�yZ��S��Ya�-{�ʇ�s? 	iF?�>���i��ۊ͕��cE��NE�>���i ���F�����L��LF��x�E}x:��j+�2���u���O���YM�HC������k J!���2������L�m
/JQ�6M4=��G�Y��a/\��cAmb_�J�9���?%�Q���r��%���G�O�֭�˴�^
�X��W�x�L��ߨVpV�ָk��٣TbqI 3�&S�(0C)W��s�ݎ�{B�"��]㮙�����~��w�%�&K0c����i �T�r{�,1�5W�5-<�:9(�H�*bBj�m̻sw��
;����;�&.��űɾ.k��ʅU�	�˒�_�3lY�c�ї���.�,n�2w%<�J'�q�Ҽ�_*2�ҵ����a����It˜[>�Ad��l��e�I���S���*�j���%�e��T��Eǳ��Z_��+~o�0K�.�GjM�no�qx��<�������Au��]�mu'��RR�p-]~j���`	��V�	*��m��,<���uC��Ӿ���M�
}f	�>���K�'�F�a�z��A��>Ē�*�c���D�ڊ���{o<F�5Ϛ`���D�+7\DA���.������oֲ���GuU��X6#��n^RF��D��hg�L�j�!��ւ��y8`~Y�5P�Vb�`	מ���ZlW�����,@����*t����