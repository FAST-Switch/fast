// megafunction wizard: %ALTLVDS%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altlvds_tx 

// ============================================================
// File Name: altera_tse_pma_lvds_tx.v
// Megafunction Name(s):
// 			altlvds_tx
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 7.2 Internal Build 97 06/25/2007 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2007 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module altera_tse_pma_lvds_tx (
	tx_in,
	tx_inclock,
	tx_out);

	input	[9:0]  tx_in;
	input	  tx_inclock;
	output	[0:0]  tx_out;

	wire [0:0] sub_wire0;
	wire [0:0] tx_out = sub_wire0[0:0];

	altlvds_tx	altlvds_tx_component (
				.tx_in (tx_in),
				.tx_inclock (tx_inclock),
				.tx_out (sub_wire0),
				.pll_areset (1'b0),
				.sync_inclock (1'b0),
				.tx_coreclock (),
				.tx_enable (1'b1),
				.tx_locked (),
				.tx_outclock (),
				.tx_pll_enable (1'b1),
				.tx_syncclock (1'b0));
	defparam
		altlvds_tx_component.common_rx_tx_pll = "ON",
		altlvds_tx_component.deserialization_factor = 10,
		altlvds_tx_component.implement_in_les = "OFF",
		altlvds_tx_component.inclock_data_alignment = "UNUSED",
		altlvds_tx_component.inclock_period = 8000,
		altlvds_tx_component.inclock_phase_shift = 0,
		altlvds_tx_component.intended_device_family = "Stratix III",
		altlvds_tx_component.lpm_type = "altlvds_tx",
		altlvds_tx_component.number_of_channels = 1,
		altlvds_tx_component.outclock_resource = "AUTO",
		altlvds_tx_component.output_data_rate = 1250,
		altlvds_tx_component.registered_input = "TX_CLKIN",
		altlvds_tx_component.use_external_pll = "OFF";


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: Clock_Choices STRING "TX_CLKIN"
// Retrieval info: PRIVATE: Clock_Mode NUMERIC "0"
// Retrieval info: PRIVATE: Data_rate STRING "1250"
// Retrieval info: PRIVATE: Deser_Factor NUMERIC "10"
// Retrieval info: PRIVATE: Enable_DPA_Mode STRING "OFF"
// Retrieval info: PRIVATE: Ext_PLL STRING "OFF"
// Retrieval info: PRIVATE: INCLOCK_PHASE_SHIFT STRING "0.00"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix III"
// Retrieval info: PRIVATE: Int_Device STRING "Stratix III"
// Retrieval info: PRIVATE: LVDS_Mode NUMERIC "0"
// Retrieval info: PRIVATE: Le_Serdes STRING "OFF"
// Retrieval info: PRIVATE: Num_Channel NUMERIC "1"
// Retrieval info: PRIVATE: OUTCLOCK_PHASE_SHIFT STRING "0.00"
// Retrieval info: PRIVATE: Outclock_Divide_By NUMERIC "10"
// Retrieval info: PRIVATE: PLL_Enable NUMERIC "0"
// Retrieval info: PRIVATE: PLL_Freq STRING "125.00"
// Retrieval info: PRIVATE: PLL_Period STRING "8.000"
// Retrieval info: PRIVATE: Reg_InOut NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: Use_Clock_Resc STRING "AUTO"
// Retrieval info: PRIVATE: Use_Common_Rx_Tx_Plls NUMERIC "1"
// Retrieval info: PRIVATE: Use_CoreClock NUMERIC "0"
// Retrieval info: PRIVATE: Use_Lock NUMERIC "0"
// Retrieval info: PRIVATE: Use_Pll_Areset NUMERIC "0"
// Retrieval info: PRIVATE: Use_Tx_Out_Phase NUMERIC "1"
// Retrieval info: CONSTANT: COMMON_RX_TX_PLL STRING "ON"
// Retrieval info: CONSTANT: DESERIALIZATION_FACTOR NUMERIC "10"
// Retrieval info: CONSTANT: IMPLEMENT_IN_LES STRING "OFF"
// Retrieval info: CONSTANT: INCLOCK_DATA_ALIGNMENT STRING "UNUSED"
// Retrieval info: CONSTANT: INCLOCK_PERIOD NUMERIC "8000"
// Retrieval info: CONSTANT: INCLOCK_PHASE_SHIFT NUMERIC "0"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix III"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altlvds_tx"
// Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "1"
// Retrieval info: CONSTANT: OUTCLOCK_RESOURCE STRING "AUTO"
// Retrieval info: CONSTANT: OUTPUT_DATA_RATE NUMERIC "1250"
// Retrieval info: CONSTANT: REGISTERED_INPUT STRING "TX_CLKIN"
// Retrieval info: CONSTANT: USE_EXTERNAL_PLL STRING "OFF"
// Retrieval info: USED_PORT: tx_in 0 0 10 0 INPUT NODEFVAL tx_in[9..0]
// Retrieval info: USED_PORT: tx_inclock 0 0 0 0 INPUT_CLK_EXT GND tx_inclock
// Retrieval info: USED_PORT: tx_out 0 0 1 0 OUTPUT NODEFVAL tx_out[0..0]
// Retrieval info: CONNECT: @tx_in 0 0 10 0 tx_in 0 0 10 0
// Retrieval info: CONNECT: tx_out 0 0 1 0 @tx_out 0 0 1 0
// Retrieval info: CONNECT: @tx_inclock 0 0 0 0 tx_inclock 0 0 0 0
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL tse_pma_lvds_tx.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL tse_pma_lvds_tx.ppf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL tse_pma_lvds_tx.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL tse_pma_lvds_tx.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL tse_pma_lvds_tx.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL tse_pma_lvds_tx_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL tse_pma_lvds_tx_bb.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_tse_pma_lvds_tx.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_tse_pma_lvds_tx.ppf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_tse_pma_lvds_tx.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_tse_pma_lvds_tx.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_tse_pma_lvds_tx.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_tse_pma_lvds_tx_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL altera_tse_pma_lvds_tx_bb.v FALSE
// Retrieval info: LIB_FILE: altera_mf
