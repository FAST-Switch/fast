��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��6�L�h�p@�
�D�i�����[�B$�N-ɛ#R \h��/6)��nJ�z)g~�HZE�x��{R6���-���r���)n�vl�ɒ-�)E��ww85��� ��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��� o�tL��nàZ�m�E*��ZQW��v�#�ͻ��n� T46��н����w�89�#�u��tJ.���Q�9���q�X��Z�(��������������Η������n���j)E�i�P�\Gj�f�Dκ�9�d��k.��-�s�+F`�9r?�4L�a�l�&�o�tƨoz�<��T����[����w���}�M�r�{���GH�����Σ��	��%�� ,a�Ew���m���8�n�7�Kr��V�I�>0ڦ<��̇���v9�_�M���}	��!r��څUѤ�<&kW���q�D�\d�+yg��32D�w�^��8��A���5�q�����e'yX�N�/T]��ن�O?�䩇h��"٭�V_q��m�ʻ-�LR�����y��ϡ#�Қ���9������M��SS�
����rO$&�^�T��AVV:�N�Ԧ��儥5s�ph����&�,� �U�}���s+i� �ҝ����'ƀ�lp�� .��&���M�r�0\R"̢���Aqb.N}.>�$Z��'͎� �UP=}q�p�����sKF��y^r
W+�;�J�ǯiz�������
�ӰS�ݚ9��0��;����E�UL?��M�C��dw��8H�M��l�r}�G]P�g>K:^a/[��h#��k�:�������T:�y�.�v���z�C�J�]M"K�*Z_����}��wm���jk���6y����F�u/��-Y��ޓ���_���`/x���%�u8'=��фԒ
��F��^|�z��X��������rw�z�{
5��w�_st��x�$}�f�#D���+��E��[�׌c%~=E���Gʡ+�2�� ��I�.��j}�!���O;��s˟��k�p^��`"��hU݆�-�@"B��#�z��:�
�|�j�*)���4i&\��9��:�yb2	��NT�b"�U�<�K�9\`�X��-_�Aj���:lSt$6���1��ol��=S�Z�Z�ψ;3}Z��e��̐ˬԖQN���-ߧ	H�$�f)�@u>n�ny���{}<f|#@@�e��q-n.���얛��]�g%�ȍ}Lg�0�֪���]q�O��\�'Ln�(C���x���i�8Q�u��\/��k|�C����[�ٹ�5�R5]�b���>b%R�y�AE�H���ȴ��D���/>� |�h�-�\�az~����^�M�z|�^>/��៎Z��O�����P'�_4����j�C�RN��5C���恄�ݕ���Bң�^���ę�����e��aN���8���z�ǋ&:/�w�H�,�Դ�q�Wu����W�#ԣ��v���gz�B�?ػ�����az�՛Zw����c_����$��bX+p)�m��-��"\�V)��[�� 0>��"p�ݛ� ��N.F/��
ۋ2��_< �0ٔOh�;��+�㲅����P��b8<��kxTob,Ք���HxZ��2��bүG����.�V
Ho���wi���������˅����3������vtp}��x��A	[p|����o�Q>��j���D�-���-��}��,��h��I�=A:-0m�i�PR�f{
�z��ae�>��0�J,�� 1��#�orz4v���~pzÎ�=�� O~���-=���Ts��q�$�<yl��޽2H��6�LE�V4+�w�1n�BN£z�\�)��A�rV8���C�3��J��Y���u���HEC}�}A�59�(��'��ud���<��k�b��Y6#ޮ���R�h�-�5]w��""Ȱ}.u��3�Q�P��ǚ�=�T;�P{�IF�8R6Vs[��	�p�I���EF�6n Q;Od�f�N���=���߫� ��pwҟ�8�0�j����T�ѽ$=��p��e��9�k-�}�����0�noZ����i�\0dE�fֿ�}���f��f"��r�<��r�%��7��]���,,8����<��\�+�.kߥ�
�_A�&xHð�ᬿ��E� �׊�`��[��L�=�K�:��1�@Xv�*+�вC̉Yo��@+TG���l9 q�����1w"U�P2������P��M�(u�*`��`	��<aS��ڭ�\�=�Y�`�������/Z��N�{Pc�0Qj~k��բ8 ��򬘰(>Q�����Z����˾r�D:�Z��tn�Ђ�y�{��m�z@�R�����C�
�= m��	pA}_C�Kћ��o����S2�'F��.´����"+;�6"�o:{�0���ػ��$���#˼|�l]t޲�;��9M����ӂ<���8�"�z����z�(Y���c�����p�W�0}�f.c[¢��+�\��D|i�:���V�O|����]�0Ff?��H@�>�т�c����at�xb8��S?�F�]nK��;rzX,�&hS�Z���kIg�o�1U��Ų�4�)��� ��o�R�v�D6�>K��Z�'z��0'g�Q}3\)���=�mJ�N��~ڔl<�D��;�|�;D�9`-E�o����+����/p^��,��*O�����[;���T:4�[v�G�ͻg�#e.���m����I?b���B��v�:�({H�$����PM�ET���4���^��H��(={r�ܨ��D�wN��8A�3H |���)��^V3��[��̊���'���v�s�K}1#��A��1r$�j0���y�^sY)	��l0���R������{	F
E���P�o�1�J�/�����!t�S@�x�}�g��	���؎1r�=��g;��M3p�8#�C)����i��AO�%fq|��%�K'��?��Uni�ۡtK�09�F�B�U�� ��B-p�5�G�ݎe�/O�B�BPd�*P7���L�*p�avx��bʩr�(�i����Ӳp�9*ƪk�f�h5R<[s��M�G!$@&V��Ik��`�s@D��fx�ؙ�G^�~q�}�p0����ܭ�25lN ��BԶE�03��<7c�W)?S�%H�a�6�n���E����S�-��czZ���	��k�8�Vc%#'B��A� ޿�qI\;�yt�nE4�q���jc�2g�OF�(@����#�J�|���JU��%*�n��&�e�(���'E&Z� �k#&1Wz9�EAb� ̸ ���G�>-߈�t+�N `�T`�s�C��n�񢱷��U[6�łq�V$a�8'dl+ !�����&��w�����Dc��)��-���t�_\4�L7$x�떃dP�,m�Ҷ�e4됉'�P���p�;�c�KѲ��v��9�Ĭ\�.�VtȾ�隃b8l�{�ҖA
q[�m�Rk�hS��<�$	����
�\�^�n'�q�{�&��K~n��P�)z��B�ڭ>����8���F��yv�5�Jg�dύÀ~<�F��t�rH�pa]��x���T������.f���q�=�X!b*����7m I�f����`��ΆWl-����y��+�	�Ϡ���ݛ2��Y� ՛,

�{�Į��
Ͼ9��;#�-b�=��\[+P��kp.| nV&��%�I�ݏ�*���%!��A��QlqW�!��\Z
;��T�z.���ά�����͚�z�m$W"yRu}��z������؋RWO"��ⷌ�x3U��Z)�e�v)�\f�H���v�Մ�8��D���#�U�1�X�(��JM���><���	/�<<JO]n`{��I�aR���]�A<�)`����A����� �ụ݅Q�|7!�X�uWC���[37HU���nY��`�ʲ�+��h��?(�� 	0^�&�^H#��w{���O�"������bC��\D�bm�:�}�71�Ԛ\8��a��d��ϝ��"ޘ�vl�ڑ>����f,��a��Iv_��?���MW9�@L���"���
.�«���Fx���O��%�1?�Ycwao��oSRPD������&����*�6�x&]�n�s�+a�e��*�i'�f��{�lC���,��^y�����-�yDf��lh�ٓ�o�	�ˎ����s�d,�=����C�ǴO���ZO�;C�� ��y�p��M�7�P5�����(�%�	G��u�Z�+|�-
d��g�?�GW��=*�)V{KX�� ����ƌ��|JsE(��l�����2�Ĭ�4����˧�qBø(� �T|N'��#=^��X9 3��ů��!qoȩ9EW��[����0��}j�+������U�՛:s��6��/��^R�bD�%.����-1J��央]��qKIMر_�y����5\�[n����(D`�'C�
�C�&�{��m̙TNr�Ɩu����p��`�1/��ýK^��G�D}�Go̤@j��k��lӰ֩M�3B��V��hd���z+��uM�=D���3YM<S2��՛irțV]�c�<o�C/a�?0~7�twZY��*��X����p�~i��6�T� ��r���w�Wkd#B��E������؟�Tz����SϳǞl^�9�Y-���-�B�#�Z0� X��H3y���܂\g�-kE�u���?����$�T��$��f���ߊ��i �=�j^��Bz�'�~O���ފk�g��o�����mT�5���
� _�+?&c[j~V��3��N��̶X>&�xN+1QM��zY�.Fon�iX�L,�:�uܦ0fql~Ť8�u�rT�1J���`/�i�c���k��%U"8��-0�݃�d���iB(��J-��	�ۋ��:zf�,3�G��\���O;���r4�Iq9�M���_�\���Y����v���`w�#3��!n-) ��8v�!Px`�9�7�F��r�����٪p圛�ֱ�=}e����s�%�ĝC� 8��&�W�P0 ./��3��A��Z]�<�;�!@�;�F**��~>�$�N� ,4�ূ� �O�LY"4>n�A�\�]��yf�/����]K,�0D�\ߚq��F����>�Ntxe����w�]� ����M�t��2m��� t'-�����Dŷ�9Ow��o���e�Y=G�{C�N�Vp�m���(� Ϊ����^r�y߲Mk.����`�*�b���J���*;Ʒ��cܵmn�@�F�iRO���8�hs�Nv�{��ӘI�o��#lj�� �����Ѓ�MP�u��+��$��
�wZ�u��CI�����v�dr+r3���B�?�f�T�:oF�}w��X�6��ˍ�F@R�A~�	�^�+?�*Q?�'�r@���'��ܹ���֞aD����)A�e��?�,�����`y(O���֎kc�n�xK��G�c,�����n�WŊˋ -3��ع�Fv?�_f�	��'s�����A�t_�2���e�i�͗���V}����ps3���t�{��1�=��=����󓜚b��:6��#{2rU3�i>�>r�